
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity CPU is
    Port ( op : in  STD_LOGIC_VECTOR (1 downto 0);
           op3 : in  STD_LOGIC_VECTOR (5 downto 0);
           salida : out  STD_LOGIC_VECTOR (5 downto 0));
end CPU;

architecture Behavioral of CPU is

begin


end Behavioral;

